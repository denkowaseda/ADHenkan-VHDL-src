library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;


entity NLAD is
     port( ADIN: in  std_logic_vector( 11 downto 0 );
           NLADOUT: out std_logic_vector( 7 downto 0 ));
end NLAD;


architecture RTL of NLAD is

signal ADIN_9 : std_logic_vector( 8 downto 0 );


begin

ADIN_9 <= ADIN(10 downto 2);

process(ADIN_9) begin

case ADIN_9 is
        when "000000000" => NLADOUT  <= "00000000" ;
        when "000000001" => NLADOUT  <= "00000111" ;
        when "000000010" => NLADOUT  <= "00001100" ;
        when "000000011" => NLADOUT  <= "00010000" ;
        when "000000100" => NLADOUT  <= "00011001" ;
        when "000000101" => NLADOUT  <= "00011100" ;
        when "000000110" => NLADOUT  <= "00011111" ;
        when "000000111" => NLADOUT  <= "00100000" ;
        when "000001000" => NLADOUT  <= "00100101" ;
        when "000001001" => NLADOUT  <= "00100111" ;
        when "000001010" => NLADOUT  <= "00101001" ;
        when "000001011" => NLADOUT  <= "00101011" ;
        when "000001100" => NLADOUT  <= "00101100" ;
        when "000001101" => NLADOUT  <= "00101110" ;
        when "000001110" => NLADOUT  <= "00101111" ;
        when "000001111" => NLADOUT  <= "00110000" ;
        when "000010000" => NLADOUT  <= "00110010" ;
        when "000010001" => NLADOUT  <= "00110011" ;
        when "000010010" => NLADOUT  <= "00110101" ;
        when "000010011" => NLADOUT  <= "00110110" ;
        when "000010100" => NLADOUT  <= "00110111" ;
        when "000010101" => NLADOUT  <= "00111000" ;
        when "000010110" => NLADOUT  <= "00111001" ;
        when "000010111" => NLADOUT  <= "00111010" ;
        when "000011000" => NLADOUT  <= "00111011" ;
        when "000011001" => NLADOUT  <= "00111100" ;
        when "000011010" => NLADOUT  <= "00111100" ;
        when "000011011" => NLADOUT  <= "00111101" ;
        when "000011100" => NLADOUT  <= "00111110" ;
        when "000011101" => NLADOUT  <= "00111111" ;
        when "000011110" => NLADOUT  <= "00111111" ;
        when "000011111" => NLADOUT  <= "01000000" ;
        when "000100000" => NLADOUT  <= "01000001" ;
        when "000100001" => NLADOUT  <= "01000001" ;
        when "000100010" => NLADOUT  <= "01000010" ;
        when "000100011" => NLADOUT  <= "01000011" ;
        when "000100100" => NLADOUT  <= "01000011" ;
        when "000100101" => NLADOUT  <= "01000100" ;
        when "000100110" => NLADOUT  <= "01000101" ;
        when "000100111" => NLADOUT  <= "01000101" ;
        when "000101000" => NLADOUT  <= "01000110" ;
        when "000101001" => NLADOUT  <= "01000110" ;
        when "000101010" => NLADOUT  <= "01000111" ;
        when "000101011" => NLADOUT  <= "01000111" ;
        when "000101100" => NLADOUT  <= "01001000" ;
        when "000101101" => NLADOUT  <= "01001000" ;
        when "000101110" => NLADOUT  <= "01001001" ;
        when "000101111" => NLADOUT  <= "01001001" ;
        when "000110000" => NLADOUT  <= "01001010" ;
        when "000110001" => NLADOUT  <= "01001010" ;
        when "000110010" => NLADOUT  <= "01001011" ;
        when "000110011" => NLADOUT  <= "01001011" ;
        when "000110100" => NLADOUT  <= "01001011" ;
        when "000110101" => NLADOUT  <= "01001100" ;
        when "000110110" => NLADOUT  <= "01001100" ;
        when "000110111" => NLADOUT  <= "01001101" ;
        when "000111000" => NLADOUT  <= "01001101" ;
        when "000111001" => NLADOUT  <= "01001110" ;
        when "000111010" => NLADOUT  <= "01001110" ;
        when "000111011" => NLADOUT  <= "01001110" ;
        when "000111100" => NLADOUT  <= "01001111" ;
        when "000111101" => NLADOUT  <= "01001111" ;
        when "000111110" => NLADOUT  <= "01001111" ;
        when "000111111" => NLADOUT  <= "01010000" ;
        when "001000000" => NLADOUT  <= "01010000" ;
        when "001000001" => NLADOUT  <= "01010000" ;
        when "001000010" => NLADOUT  <= "01010001" ;
        when "001000011" => NLADOUT  <= "01010001" ;
        when "001000100" => NLADOUT  <= "01010001" ;
        when "001000101" => NLADOUT  <= "01010010" ;
        when "001000110" => NLADOUT  <= "01010010" ;
        when "001000111" => NLADOUT  <= "01010010" ;
        when "001001000" => NLADOUT  <= "01010011" ;
        when "001001001" => NLADOUT  <= "01010011" ;
        when "001001010" => NLADOUT  <= "01010011" ;
        when "001001011" => NLADOUT  <= "01010100" ;
        when "001001100" => NLADOUT  <= "01010100" ;
        when "001001101" => NLADOUT  <= "01010100" ;
        when "001001110" => NLADOUT  <= "01010101" ;
        when "001001111" => NLADOUT  <= "01010101" ;
        when "001010000" => NLADOUT  <= "01010101" ;
        when "001010001" => NLADOUT  <= "01010101" ;
        when "001010010" => NLADOUT  <= "01010110" ;
        when "001010011" => NLADOUT  <= "01010110" ;
        when "001010100" => NLADOUT  <= "01010110" ;
        when "001010101" => NLADOUT  <= "01010110" ;
        when "001010110" => NLADOUT  <= "01010111" ;
        when "001010111" => NLADOUT  <= "01010111" ;
        when "001011000" => NLADOUT  <= "01010111" ;
        when "001011001" => NLADOUT  <= "01011000" ;
        when "001011010" => NLADOUT  <= "01011000" ;
        when "001011011" => NLADOUT  <= "01011000" ;
        when "001011100" => NLADOUT  <= "01011000" ;
        when "001011101" => NLADOUT  <= "01011001" ;
        when "001011110" => NLADOUT  <= "01011001" ;
        when "001011111" => NLADOUT  <= "01011001" ;
        when "001100000" => NLADOUT  <= "01011001" ;
        when "001100001" => NLADOUT  <= "01011001" ;
        when "001100010" => NLADOUT  <= "01011010" ;
        when "001100011" => NLADOUT  <= "01011010" ;
        when "001100100" => NLADOUT  <= "01011010" ;
        when "001100101" => NLADOUT  <= "01011010" ;
        when "001100110" => NLADOUT  <= "01011011" ;
        when "001100111" => NLADOUT  <= "01011011" ;
        when "001101000" => NLADOUT  <= "01011011" ;
        when "001101001" => NLADOUT  <= "01011011" ;
        when "001101010" => NLADOUT  <= "01011011" ;
        when "001101011" => NLADOUT  <= "01011100" ;
        when "001101100" => NLADOUT  <= "01011100" ;
        when "001101101" => NLADOUT  <= "01011100" ;
        when "001101110" => NLADOUT  <= "01011100" ;
        when "001101111" => NLADOUT  <= "01011101" ;
        when "001110000" => NLADOUT  <= "01011101" ;
        when "001110001" => NLADOUT  <= "01011101" ;
        when "001110010" => NLADOUT  <= "01011101" ;
        when "001110011" => NLADOUT  <= "01011101" ;
        when "001110100" => NLADOUT  <= "01011110" ;
        when "001110101" => NLADOUT  <= "01011110" ;
        when "001110110" => NLADOUT  <= "01011110" ;
        when "001110111" => NLADOUT  <= "01011110" ;
        when "001111000" => NLADOUT  <= "01011110" ;
        when "001111001" => NLADOUT  <= "01011110" ;
        when "001111010" => NLADOUT  <= "01011111" ;
        when "001111011" => NLADOUT  <= "01011111" ;
        when "001111100" => NLADOUT  <= "01011111" ;
        when "001111101" => NLADOUT  <= "01011111" ;
        when "001111110" => NLADOUT  <= "01011111" ;
        when "001111111" => NLADOUT  <= "01100000" ;
        when "010000000" => NLADOUT  <= "01100000" ;
        when "010000001" => NLADOUT  <= "01100000" ;
        when "010000010" => NLADOUT  <= "01100000" ;
        when "010000011" => NLADOUT  <= "01100000" ;
        when "010000100" => NLADOUT  <= "01100000" ;
        when "010000101" => NLADOUT  <= "01100001" ;
        when "010000110" => NLADOUT  <= "01100001" ;
        when "010000111" => NLADOUT  <= "01100001" ;
        when "010001000" => NLADOUT  <= "01100001" ;
        when "010001001" => NLADOUT  <= "01100001" ;
        when "010001010" => NLADOUT  <= "01100001" ;
        when "010001011" => NLADOUT  <= "01100010" ;
        when "010001100" => NLADOUT  <= "01100010" ;
        when "010001101" => NLADOUT  <= "01100010" ;
        when "010001110" => NLADOUT  <= "01100010" ;
        when "010001111" => NLADOUT  <= "01100010" ;
        when "010010000" => NLADOUT  <= "01100010" ;
        when "010010001" => NLADOUT  <= "01100011" ;
        when "010010010" => NLADOUT  <= "01100011" ;
        when "010010011" => NLADOUT  <= "01100011" ;
        when "010010100" => NLADOUT  <= "01100011" ;
        when "010010101" => NLADOUT  <= "01100011" ;
        when "010010110" => NLADOUT  <= "01100011" ;
        when "010010111" => NLADOUT  <= "01100100" ;
        when "010011000" => NLADOUT  <= "01100100" ;
        when "010011001" => NLADOUT  <= "01100100" ;
        when "010011010" => NLADOUT  <= "01100100" ;
        when "010011011" => NLADOUT  <= "01100100" ;
        when "010011100" => NLADOUT  <= "01100100" ;
        when "010011101" => NLADOUT  <= "01100100" ;
        when "010011110" => NLADOUT  <= "01100101" ;
        when "010011111" => NLADOUT  <= "01100101" ;
        when "010100000" => NLADOUT  <= "01100101" ;
        when "010100001" => NLADOUT  <= "01100101" ;
        when "010100010" => NLADOUT  <= "01100101" ;
        when "010100011" => NLADOUT  <= "01100101" ;
        when "010100100" => NLADOUT  <= "01100101" ;
        when "010100101" => NLADOUT  <= "01100110" ;
        when "010100110" => NLADOUT  <= "01100110" ;
        when "010100111" => NLADOUT  <= "01100110" ;
        when "010101000" => NLADOUT  <= "01100110" ;
        when "010101001" => NLADOUT  <= "01100110" ;
        when "010101010" => NLADOUT  <= "01100110" ;
        when "010101011" => NLADOUT  <= "01100110" ;
        when "010101100" => NLADOUT  <= "01100110" ;
        when "010101101" => NLADOUT  <= "01100111" ;
        when "010101110" => NLADOUT  <= "01100111" ;
        when "010101111" => NLADOUT  <= "01100111" ;
        when "010110000" => NLADOUT  <= "01100111" ;
        when "010110001" => NLADOUT  <= "01100111" ;
        when "010110010" => NLADOUT  <= "01100111" ;
        when "010110011" => NLADOUT  <= "01100111" ;
        when "010110100" => NLADOUT  <= "01101000" ;
        when "010110101" => NLADOUT  <= "01101000" ;
        when "010110110" => NLADOUT  <= "01101000" ;
        when "010110111" => NLADOUT  <= "01101000" ;
        when "010111000" => NLADOUT  <= "01101000" ;
        when "010111001" => NLADOUT  <= "01101000" ;
        when "010111010" => NLADOUT  <= "01101000" ;
        when "010111011" => NLADOUT  <= "01101000" ;
        when "010111100" => NLADOUT  <= "01101001" ;
        when "010111101" => NLADOUT  <= "01101001" ;
        when "010111110" => NLADOUT  <= "01101001" ;
        when "010111111" => NLADOUT  <= "01101001" ;
        when "011000000" => NLADOUT  <= "01101001" ;
        when "011000001" => NLADOUT  <= "01101001" ;
        when "011000010" => NLADOUT  <= "01101001" ;
        when "011000011" => NLADOUT  <= "01101001" ;
        when "011000100" => NLADOUT  <= "01101001" ;
        when "011000101" => NLADOUT  <= "01101010" ;
        when "011000110" => NLADOUT  <= "01101010" ;
        when "011000111" => NLADOUT  <= "01101010" ;
        when "011001000" => NLADOUT  <= "01101010" ;
        when "011001001" => NLADOUT  <= "01101010" ;
        when "011001010" => NLADOUT  <= "01101010" ;
        when "011001011" => NLADOUT  <= "01101010" ;
        when "011001100" => NLADOUT  <= "01101010" ;
        when "011001101" => NLADOUT  <= "01101010" ;
        when "011001110" => NLADOUT  <= "01101011" ;
        when "011001111" => NLADOUT  <= "01101011" ;
        when "011010000" => NLADOUT  <= "01101011" ;
        when "011010001" => NLADOUT  <= "01101011" ;
        when "011010010" => NLADOUT  <= "01101011" ;
        when "011010011" => NLADOUT  <= "01101011" ;
        when "011010100" => NLADOUT  <= "01101011" ;
        when "011010101" => NLADOUT  <= "01101011" ;
        when "011010110" => NLADOUT  <= "01101011" ;
        when "011010111" => NLADOUT  <= "01101100" ;
        when "011011000" => NLADOUT  <= "01101100" ;
        when "011011001" => NLADOUT  <= "01101100" ;
        when "011011010" => NLADOUT  <= "01101100" ;
        when "011011011" => NLADOUT  <= "01101100" ;
        when "011011100" => NLADOUT  <= "01101100" ;
        when "011011101" => NLADOUT  <= "01101100" ;
        when "011011110" => NLADOUT  <= "01101100" ;
        when "011011111" => NLADOUT  <= "01101100" ;
        when "011100000" => NLADOUT  <= "01101101" ;
        when "011100001" => NLADOUT  <= "01101101" ;
        when "011100010" => NLADOUT  <= "01101101" ;
        when "011100011" => NLADOUT  <= "01101101" ;
        when "011100100" => NLADOUT  <= "01101101" ;
        when "011100101" => NLADOUT  <= "01101101" ;
        when "011100110" => NLADOUT  <= "01101101" ;
        when "011100111" => NLADOUT  <= "01101101" ;
        when "011101000" => NLADOUT  <= "01101101" ;
        when "011101001" => NLADOUT  <= "01101101" ;
        when "011101010" => NLADOUT  <= "01101110" ;
        when "011101011" => NLADOUT  <= "01101110" ;
        when "011101100" => NLADOUT  <= "01101110" ;
        when "011101101" => NLADOUT  <= "01101110" ;
        when "011101110" => NLADOUT  <= "01101110" ;
        when "011101111" => NLADOUT  <= "01101110" ;
        when "011110000" => NLADOUT  <= "01101110" ;
        when "011110001" => NLADOUT  <= "01101110" ;
        when "011110010" => NLADOUT  <= "01101110" ;
        when "011110011" => NLADOUT  <= "01101110" ;
        when "011110100" => NLADOUT  <= "01101110" ;
        when "011110101" => NLADOUT  <= "01101111" ;
        when "011110110" => NLADOUT  <= "01101111" ;
        when "011110111" => NLADOUT  <= "01101111" ;
        when "011111000" => NLADOUT  <= "01101111" ;
        when "011111001" => NLADOUT  <= "01101111" ;
        when "011111010" => NLADOUT  <= "01101111" ;
        when "011111011" => NLADOUT  <= "01101111" ;
        when "011111100" => NLADOUT  <= "01101111" ;
        when "011111101" => NLADOUT  <= "01101111" ;
        when "011111110" => NLADOUT  <= "01101111" ;
        when "011111111" => NLADOUT  <= "01101111" ;
        when "100000000" => NLADOUT  <= "01110000" ;
        when "100000001" => NLADOUT  <= "01110000" ;
        when "100000010" => NLADOUT  <= "01110000" ;
        when "100000011" => NLADOUT  <= "01110000" ;
        when "100000100" => NLADOUT  <= "01110000" ;
        when "100000101" => NLADOUT  <= "01110000" ;
        when "100000110" => NLADOUT  <= "01110000" ;
        when "100000111" => NLADOUT  <= "01110000" ;
        when "100001000" => NLADOUT  <= "01110000" ;
        when "100001001" => NLADOUT  <= "01110000" ;
        when "100001010" => NLADOUT  <= "01110000" ;
        when "100001011" => NLADOUT  <= "01110001" ;
        when "100001100" => NLADOUT  <= "01110001" ;
        when "100001101" => NLADOUT  <= "01110001" ;
        when "100001110" => NLADOUT  <= "01110001" ;
        when "100001111" => NLADOUT  <= "01110001" ;
        when "100010000" => NLADOUT  <= "01110001" ;
        when "100010001" => NLADOUT  <= "01110001" ;
        when "100010010" => NLADOUT  <= "01110001" ;
        when "100010011" => NLADOUT  <= "01110001" ;
        when "100010100" => NLADOUT  <= "01110001" ;
        when "100010101" => NLADOUT  <= "01110001" ;
        when "100010110" => NLADOUT  <= "01110001" ;
        when "100010111" => NLADOUT  <= "01110010" ;
        when "100011000" => NLADOUT  <= "01110010" ;
        when "100011001" => NLADOUT  <= "01110010" ;
        when "100011010" => NLADOUT  <= "01110010" ;
        when "100011011" => NLADOUT  <= "01110010" ;
        when "100011100" => NLADOUT  <= "01110010" ;
        when "100011101" => NLADOUT  <= "01110010" ;
        when "100011110" => NLADOUT  <= "01110010" ;
        when "100011111" => NLADOUT  <= "01110010" ;
        when "100100000" => NLADOUT  <= "01110010" ;
        when "100100001" => NLADOUT  <= "01110010" ;
        when "100100010" => NLADOUT  <= "01110010" ;
        when "100100011" => NLADOUT  <= "01110011" ;
        when "100100100" => NLADOUT  <= "01110011" ;
        when "100100101" => NLADOUT  <= "01110011" ;
        when "100100110" => NLADOUT  <= "01110011" ;
        when "100100111" => NLADOUT  <= "01110011" ;
        when "100101000" => NLADOUT  <= "01110011" ;
        when "100101001" => NLADOUT  <= "01110011" ;
        when "100101010" => NLADOUT  <= "01110011" ;
        when "100101011" => NLADOUT  <= "01110011" ;
        when "100101100" => NLADOUT  <= "01110011" ;
        when "100101101" => NLADOUT  <= "01110011" ;
        when "100101110" => NLADOUT  <= "01110011" ;
        when "100101111" => NLADOUT  <= "01110011" ;
        when "100110000" => NLADOUT  <= "01110100" ;
        when "100110001" => NLADOUT  <= "01110100" ;
        when "100110010" => NLADOUT  <= "01110100" ;
        when "100110011" => NLADOUT  <= "01110100" ;
        when "100110100" => NLADOUT  <= "01110100" ;
        when "100110101" => NLADOUT  <= "01110100" ;
        when "100110110" => NLADOUT  <= "01110100" ;
        when "100110111" => NLADOUT  <= "01110100" ;
        when "100111000" => NLADOUT  <= "01110100" ;
        when "100111001" => NLADOUT  <= "01110100" ;
        when "100111010" => NLADOUT  <= "01110100" ;
        when "100111011" => NLADOUT  <= "01110100" ;
        when "100111100" => NLADOUT  <= "01110100" ;
        when "100111101" => NLADOUT  <= "01110100" ;
        when "100111110" => NLADOUT  <= "01110101" ;
        when "100111111" => NLADOUT  <= "01110101" ;
        when "101000000" => NLADOUT  <= "01110101" ;
        when "101000001" => NLADOUT  <= "01110101" ;
        when "101000010" => NLADOUT  <= "01110101" ;
        when "101000011" => NLADOUT  <= "01110101" ;
        when "101000100" => NLADOUT  <= "01110101" ;
        when "101000101" => NLADOUT  <= "01110101" ;
        when "101000110" => NLADOUT  <= "01110101" ;
        when "101000111" => NLADOUT  <= "01110101" ;
        when "101001000" => NLADOUT  <= "01110101" ;
        when "101001001" => NLADOUT  <= "01110101" ;
        when "101001010" => NLADOUT  <= "01110101" ;
        when "101001011" => NLADOUT  <= "01110101" ;
        when "101001100" => NLADOUT  <= "01110110" ;
        when "101001101" => NLADOUT  <= "01110110" ;
        when "101001110" => NLADOUT  <= "01110110" ;
        when "101001111" => NLADOUT  <= "01110110" ;
        when "101010000" => NLADOUT  <= "01110110" ;
        when "101010001" => NLADOUT  <= "01110110" ;
        when "101010010" => NLADOUT  <= "01110110" ;
        when "101010011" => NLADOUT  <= "01110110" ;
        when "101010100" => NLADOUT  <= "01110110" ;
        when "101010101" => NLADOUT  <= "01110110" ;
        when "101010110" => NLADOUT  <= "01110110" ;
        when "101010111" => NLADOUT  <= "01110110" ;
        when "101011000" => NLADOUT  <= "01110110" ;
        when "101011001" => NLADOUT  <= "01110110" ;
        when "101011010" => NLADOUT  <= "01110110" ;
        when "101011011" => NLADOUT  <= "01110111" ;
        when "101011100" => NLADOUT  <= "01110111" ;
        when "101011101" => NLADOUT  <= "01110111" ;
        when "101011110" => NLADOUT  <= "01110111" ;
        when "101011111" => NLADOUT  <= "01110111" ;
        when "101100000" => NLADOUT  <= "01110111" ;
        when "101100001" => NLADOUT  <= "01110111" ;
        when "101100010" => NLADOUT  <= "01110111" ;
        when "101100011" => NLADOUT  <= "01110111" ;
        when "101100100" => NLADOUT  <= "01110111" ;
        when "101100101" => NLADOUT  <= "01110111" ;
        when "101100110" => NLADOUT  <= "01110111" ;
        when "101100111" => NLADOUT  <= "01110111" ;
        when "101101000" => NLADOUT  <= "01110111" ;
        when "101101001" => NLADOUT  <= "01110111" ;
        when "101101010" => NLADOUT  <= "01111000" ;
        when "101101011" => NLADOUT  <= "01111000" ;
        when "101101100" => NLADOUT  <= "01111000" ;
        when "101101101" => NLADOUT  <= "01111000" ;
        when "101101110" => NLADOUT  <= "01111000" ;
        when "101101111" => NLADOUT  <= "01111000" ;
        when "101110000" => NLADOUT  <= "01111000" ;
        when "101110001" => NLADOUT  <= "01111000" ;
        when "101110010" => NLADOUT  <= "01111000" ;
        when "101110011" => NLADOUT  <= "01111000" ;
        when "101110100" => NLADOUT  <= "01111000" ;
        when "101110101" => NLADOUT  <= "01111000" ;
        when "101110110" => NLADOUT  <= "01111000" ;
        when "101110111" => NLADOUT  <= "01111000" ;
        when "101111000" => NLADOUT  <= "01111000" ;
        when "101111001" => NLADOUT  <= "01111000" ;
        when "101111010" => NLADOUT  <= "01111001" ;
        when "101111011" => NLADOUT  <= "01111001" ;
        when "101111100" => NLADOUT  <= "01111001" ;
        when "101111101" => NLADOUT  <= "01111001" ;
        when "101111110" => NLADOUT  <= "01111001" ;
        when "101111111" => NLADOUT  <= "01111001" ;
        when "110000000" => NLADOUT  <= "01111001" ;
        when "110000001" => NLADOUT  <= "01111001" ;
        when "110000010" => NLADOUT  <= "01111001" ;
        when "110000011" => NLADOUT  <= "01111001" ;
        when "110000100" => NLADOUT  <= "01111001" ;
        when "110000101" => NLADOUT  <= "01111001" ;
        when "110000110" => NLADOUT  <= "01111001" ;
        when "110000111" => NLADOUT  <= "01111001" ;
        when "110001000" => NLADOUT  <= "01111001" ;
        when "110001001" => NLADOUT  <= "01111001" ;
        when "110001010" => NLADOUT  <= "01111001" ;
        when "110001011" => NLADOUT  <= "01111010" ;
        when "110001100" => NLADOUT  <= "01111010" ;
        when "110001101" => NLADOUT  <= "01111010" ;
        when "110001110" => NLADOUT  <= "01111010" ;
        when "110001111" => NLADOUT  <= "01111010" ;
        when "110010000" => NLADOUT  <= "01111010" ;
        when "110010001" => NLADOUT  <= "01111010" ;
        when "110010010" => NLADOUT  <= "01111010" ;
        when "110010011" => NLADOUT  <= "01111010" ;
        when "110010100" => NLADOUT  <= "01111010" ;
        when "110010101" => NLADOUT  <= "01111010" ;
        when "110010110" => NLADOUT  <= "01111010" ;
        when "110010111" => NLADOUT  <= "01111010" ;
        when "110011000" => NLADOUT  <= "01111010" ;
        when "110011001" => NLADOUT  <= "01111010" ;
        when "110011010" => NLADOUT  <= "01111010" ;
        when "110011011" => NLADOUT  <= "01111010" ;
        when "110011100" => NLADOUT  <= "01111010" ;
        when "110011101" => NLADOUT  <= "01111011" ;
        when "110011110" => NLADOUT  <= "01111011" ;
        when "110011111" => NLADOUT  <= "01111011" ;
        when "110100000" => NLADOUT  <= "01111011" ;
        when "110100001" => NLADOUT  <= "01111011" ;
        when "110100010" => NLADOUT  <= "01111011" ;
        when "110100011" => NLADOUT  <= "01111011" ;
        when "110100100" => NLADOUT  <= "01111011" ;
        when "110100101" => NLADOUT  <= "01111011" ;
        when "110100110" => NLADOUT  <= "01111011" ;
        when "110100111" => NLADOUT  <= "01111011" ;
        when "110101000" => NLADOUT  <= "01111011" ;
        when "110101001" => NLADOUT  <= "01111011" ;
        when "110101010" => NLADOUT  <= "01111011" ;
        when "110101011" => NLADOUT  <= "01111011" ;
        when "110101100" => NLADOUT  <= "01111011" ;
        when "110101101" => NLADOUT  <= "01111011" ;
        when "110101110" => NLADOUT  <= "01111011" ;
        when "110101111" => NLADOUT  <= "01111100" ;
        when "110110000" => NLADOUT  <= "01111100" ;
        when "110110001" => NLADOUT  <= "01111100" ;
        when "110110010" => NLADOUT  <= "01111100" ;
        when "110110011" => NLADOUT  <= "01111100" ;
        when "110110100" => NLADOUT  <= "01111100" ;
        when "110110101" => NLADOUT  <= "01111100" ;
        when "110110110" => NLADOUT  <= "01111100" ;
        when "110110111" => NLADOUT  <= "01111100" ;
        when "110111000" => NLADOUT  <= "01111100" ;
        when "110111001" => NLADOUT  <= "01111100" ;
        when "110111010" => NLADOUT  <= "01111100" ;
        when "110111011" => NLADOUT  <= "01111100" ;
        when "110111100" => NLADOUT  <= "01111100" ;
        when "110111101" => NLADOUT  <= "01111100" ;
        when "110111110" => NLADOUT  <= "01111100" ;
        when "110111111" => NLADOUT  <= "01111100" ;
        when "111000000" => NLADOUT  <= "01111100" ;
        when "111000001" => NLADOUT  <= "01111100" ;
        when "111000010" => NLADOUT  <= "01111101" ;
        when "111000011" => NLADOUT  <= "01111101" ;
        when "111000100" => NLADOUT  <= "01111101" ;
        when "111000101" => NLADOUT  <= "01111101" ;
        when "111000110" => NLADOUT  <= "01111101" ;
        when "111000111" => NLADOUT  <= "01111101" ;
        when "111001000" => NLADOUT  <= "01111101" ;
        when "111001001" => NLADOUT  <= "01111101" ;
        when "111001010" => NLADOUT  <= "01111101" ;
        when "111001011" => NLADOUT  <= "01111101" ;
        when "111001100" => NLADOUT  <= "01111101" ;
        when "111001101" => NLADOUT  <= "01111101" ;
        when "111001110" => NLADOUT  <= "01111101" ;
        when "111001111" => NLADOUT  <= "01111101" ;
        when "111010000" => NLADOUT  <= "01111101" ;
        when "111010001" => NLADOUT  <= "01111101" ;
        when "111010010" => NLADOUT  <= "01111101" ;
        when "111010011" => NLADOUT  <= "01111101" ;
        when "111010100" => NLADOUT  <= "01111101" ;
        when "111010101" => NLADOUT  <= "01111101" ;
        when "111010110" => NLADOUT  <= "01111110" ;
        when "111010111" => NLADOUT  <= "01111110" ;
        when "111011000" => NLADOUT  <= "01111110" ;
        when "111011001" => NLADOUT  <= "01111110" ;
        when "111011010" => NLADOUT  <= "01111110" ;
        when "111011011" => NLADOUT  <= "01111110" ;
        when "111011100" => NLADOUT  <= "01111110" ;
        when "111011101" => NLADOUT  <= "01111110" ;
        when "111011110" => NLADOUT  <= "01111110" ;
        when "111011111" => NLADOUT  <= "01111110" ;
        when "111100000" => NLADOUT  <= "01111110" ;
        when "111100001" => NLADOUT  <= "01111110" ;
        when "111100010" => NLADOUT  <= "01111110" ;
        when "111100011" => NLADOUT  <= "01111110" ;
        when "111100100" => NLADOUT  <= "01111110" ;
        when "111100101" => NLADOUT  <= "01111110" ;
        when "111100110" => NLADOUT  <= "01111110" ;
        when "111100111" => NLADOUT  <= "01111110" ;
        when "111101000" => NLADOUT  <= "01111110" ;
        when "111101001" => NLADOUT  <= "01111110" ;
        when "111101010" => NLADOUT  <= "01111110" ;
        when "111101011" => NLADOUT  <= "01111111" ;
        when "111101100" => NLADOUT  <= "01111111" ;
        when "111101101" => NLADOUT  <= "01111111" ;
        when "111101110" => NLADOUT  <= "01111111" ;
        when "111101111" => NLADOUT  <= "01111111" ;
        when "111110000" => NLADOUT  <= "01111111" ;
        when "111110001" => NLADOUT  <= "01111111" ;
        when "111110010" => NLADOUT  <= "01111111" ;
        when "111110011" => NLADOUT  <= "01111111" ;
        when "111110100" => NLADOUT  <= "01111111" ;
        when "111110101" => NLADOUT  <= "01111111" ;
        when "111110110" => NLADOUT  <= "01111111" ;
        when "111110111" => NLADOUT  <= "01111111" ;
        when "111111000" => NLADOUT  <= "01111111" ;
        when "111111001" => NLADOUT  <= "01111111" ;
        when "111111010" => NLADOUT  <= "01111111" ;
        when "111111011" => NLADOUT  <= "01111111" ;
        when "111111100" => NLADOUT  <= "01111111" ;
        when "111111101" => NLADOUT  <= "01111111" ;
        when "111111110" => NLADOUT  <= "01111111" ;
        when "111111111" => NLADOUT  <= "01111111" ;
        when  others     => NLADOUT  <= "00000000" ;
end case;

end process;

end RTL;

